module bcdmapper(
    input wire [3:0] BCD,
    output wire [7:0] segment
);

    assign segment = ((BCD == 4'b0000) ? 8'b11111100 : 8'b00000000
    | (BCD == 4'b0001) ? 8'b01100000 : 8'b00000000
    | (BCD == 4'b0010) ? 8'b11011010 : 8'b00000000
    | (BCD == 4'b0011) ? 8'b11110010 : 8'b00000000
    | (BCD == 4'b0100) ? 8'b01100110 : 8'b00000000
    | (BCD == 4'b0101) ? 8'b10110110 : 8'b00000000
    | (BCD == 4'b0110) ? 8'b10111110 : 8'b00000000
    | (BCD == 4'b0111) ? 8'b11100000 : 8'b00000000
    | (BCD == 4'b1000) ? 8'b11111110 : 8'b00000000
    | (BCD == 4'b1001) ? 8'b11110110 : 8'b00000000 // 9
    | (BCD == 4'b1010) ? 8'b11101110 : 8'b00000000 // A
    | (BCD == 4'b1011) ? 8'b00111110 : 8'b00000000
    | (BCD == 4'b1100) ? 8'b10011100 : 8'b00000000
    | (BCD == 4'b1101) ? 8'b01111010 : 8'b00000000
    | (BCD == 4'b1110) ? 8'b10011110 : 8'b00000000
    | (BCD == 4'b1111) ? 8'b10001110 : 8'b00000000);

endmodule
